// "Monitor" core that is loaded as the default core on power-up.
// nand2mario, 2025.2

`ifndef VERILATOR
`ifndef MEGA
`ifndef CONSOLE
`ifndef PRIMER
`ifndef NANO
`error "config.v must be read before monitor_top.v"
`endif
`endif
`endif
`endif
`endif

import configPackage::*;

module monitor_top (
    input        sys_clk,
    input        s0,

    // UART
    input        UART_RXD,
    output       UART_TXD,

    // HDMI TX
    output       tmds_clk_p,    
    output       tmds_clk_n,
    output [2:0] tmds_d_p,
    output [2:0] tmds_d_n,

    // USB1 and USB2
`ifdef USB1
    inout usb1_dp,
    inout usb1_dn,
`endif
`ifdef USB2
    inout usb2_dp,
    inout usb2_dn,
`endif

`ifdef CONTROLLER_SNES
    // snes controllers
    output       joy1_strb,
    output       joy1_clk,
    input        joy1_data,
    output       joy2_strb,
    output       joy2_clk,
    input        joy2_data,
`endif

`ifdef CONTROLLER_DS2
    // dualshock controllers
    output       ds_clk,
    input        ds_miso,
    output       ds_mosi,
    output       ds_cs,
    output       ds_clk2,
    input        ds_miso2,
    output       ds_mosi2,
    output       ds_cs2,
`endif

    // LED
    output [7:0] led
);

// Clock signals
wire clk;                       // main clock 50Mhz
wire clk27;                     // 27Mhz for HDMI
wire hclk5, hclk;               // 720p pixel clock at 74.25Mhz, and 5x high-speed

reg resetn = 0;              // reset is cleared after 4 cycles

// HDMI clocks
`ifdef NANO
// GW2A Nano20K
assign clk27 = sys_clk;       
assign clk = sys_clk;
localparam FREQ = 27_000_000;
gowin_pll_hdmi pll_hdmi (.clkin(clk27), .clkout(hclk5));
CLKDIV #(.DIV_MODE(5)) div5 (
    .CLKOUT(hclk),
    .HCLKIN(hclk5),
    .RESETN(1'b1),
    .CALIB(1'b0)
);

`else
// GW5 devices
assign clk = sys_clk;
localparam FREQ = 50_000_000;
pll_27 pll_27 (
    .clkin(sys_clk),
    .clkout0(clk27)
);
pll_74 pll_74 (
    .clkin(clk27),              // 27 Mhz input
    .clkout0(hclk), .clkout1(hclk5)
);
`endif

reg [15:0] resetcnt = 16'hffff;
always @(posedge clk) begin
    resetcnt <= resetcnt == 0 ? 0 : resetcnt - 1;
     if (resetcnt == 0)
//  if (resetcnt == 0 && s0)    // primer25k, nano20k
//  if (resetcnt == 0 && ~s0)   // mega138k
        resetn <= 1'b1;
end

wire overlay;
wor [11:0] joy1_btns, joy2_btns;

// Controller input
`ifdef CONTROLLER_SNES
controller_snes #(.FREQ(FREQ)) joy1_snes (
    .clk(clk), .resetn(resetn), .buttons(joy1_btns),
    .joy_strb(joy1_strb), .joy_clk(joy1_clk), .joy_data(joy1_data)
);
controller_snes #(.FREQ(FREQ)) joy2_snes (
    .clk(clk), .resetn(resetn), .buttons(joy2_btns),
    .joy_strb(joy2_strb), .joy_clk(joy2_clk), .joy_data(joy2_data)
);
`endif

`ifdef CONTROLLER_DS2
controller_ds2 #(.FREQ(FREQ)) joy1_ds2 (
    .clk(clk), .snes_buttons(joy1_btns),
    .ds_clk(ds_clk), .ds_miso(ds_miso), .ds_mosi(ds_mosi), .ds_cs(ds_cs) 
);
controller_ds2 #(.FREQ(FREQ)) joy2_ds2 (
   .clk(clk), .snes_buttons(joy2_btns),
   .ds_clk(ds_clk2), .ds_miso(ds_miso2), .ds_mosi(ds_mosi2), .ds_cs(ds_cs2) 
);
`endif

wire [11:0] joy_usb1, joy_usb2;

`ifdef USB1
wire clk12;
wire pll_lock_12;
wire usb_conerr;
wire [1:0] usb_type;
pll_12 pll12(.clkin(sys_clk), .clkout0(clk12), .lock(pll_lock_12));
usb_hid_host usb_hid_host (
    .usbclk(clk12), .usbrst_n(pll_lock_12),
    .usb_dm(usb1_dn), .usb_dp(usb1_dp),
    .game_snes(joy_usb1), .typ(usb_type), .conerr(usb_conerr)
);
assign led = ~{joy_usb1[4:0], usb_type, usb_conerr};
`else
assign joy_usb1 = 12'b0;
`endif

`ifdef USB2
usb_hid_host usb_hid_host2 (
    .usbclk(clk12), .usbrst_n(pll_lock_12),
    .usb_dm(usb2_dn), .usb_dp(usb2_dp),
    .game_snes(joy_usb2)
);
`else
assign joy_usb2 = 12'b0;
`endif

wire [14:0] overlay_color;
wire [7:0] overlay_x;
wire [7:0] overlay_y;

monitor2hdmi s2h(
    .clk(clk), .resetn(1'b1), 
    .overlay(overlay), .overlay_x(overlay_x), .overlay_y(overlay_y),
    .overlay_color(overlay_color), 
    .clk_pixel(hclk),.clk_5x_pixel(hclk5),
    .tmds_clk_n(tmds_clk_n), .tmds_clk_p(tmds_clk_p),
    .tmds_d_n(tmds_d_n), .tmds_d_p(tmds_d_p)
);

// IOSys for menu, rom loading...
iosys_bl616 #(.CORE_ID(0), .FREQ(FREQ), .COLOR_LOGO(15'b11011_10010_00011)) sys (        // CORE ID 0: Monitor
    .clk(clk), .hclk(hclk), .resetn(resetn),
    // overlay generated by textdisp
    .overlay(overlay), .overlay_x(overlay_x), .overlay_y(overlay_y), .overlay_color(overlay_color),
    // joystick buttons to be sent to companion MCU
    .joy1(joy1_btns | joy_usb1), .joy2(joy2_btns | joy_usb2),
    // UART connection to the companion MCU
    .uart_rx(UART_RXD), .uart_tx(UART_TXD)
);

endmodule
