// "Monitor" core that is loaded as the default core on power-up.
// nand2mario, 2025.2

`ifndef VERILATOR
`ifndef MEGA
`ifndef CONSOLE
`error "config.v must be read before snestang_top.v"
`endif
`endif
`endif

import configPackage::*;

module monitor_top (
    input        sys_clk,
    input        s0,

    // UART
    input        UART_RXD,
    output       UART_TXD,

    // HDMI TX
    output       tmds_clk_p,    
    output       tmds_clk_n,
    output [2:0] tmds_d_p,
    output [2:0] tmds_d_n,

    // Slave SPI to companion MCU
    input        sspi_clk;      
    input        sspi_cs;
    input        sspi_mosi;
    output       sspi_miso;

`ifdef CONTROLLER_SNES
    // snes controllers
    output       joy1_strb,
    output       joy1_clk,
    input        joy1_data,
    output       joy2_strb,
    output       joy2_clk,
    input        joy2_data,
`endif

`ifdef CONTROLLER_DS2
    // dualshock controllers
    output       ds_clk,
    input        ds_miso,
    output       ds_mosi,
    output       ds_cs,
    output       ds_clk2,
    input        ds_miso2,
    output       ds_mosi2,
    output       ds_cs2,
`endif

    // LED
    output [1:0] led
);

// Clock signals
wire clk = sys_clk;             // main clock 50Mhz
wire clk27;                     // 27Mhz for HDMI
wire hclk5, hclk;               // 720p pixel clock at 74.25Mhz, and 5x high-speed

reg resetn = 1'b0;              // reset is cleared after 4 cycles

reg [15:0] resetcnt = 16'hffff;
always @(posedge mclk) begin
    resetcnt <= resetcnt == 0 ? 0 : resetcnt - 1;
     if (resetcnt == 0)
//  if (resetcnt == 0 && s0)   // primer25k, nano20k
//     if (resetcnt == 0 && ~s0)   // mega138k
        resetn <= 1'b1;
end

// HDMI clocks
gowin_pll_27 pll_27 (
    .clkin(sys_clk),
    .clkout0(clk27)
);
gowin_pll_hdmi pll_hdmi (
    .clkin(clk27),              // 27 Mhz input
    .clkout0(hclk5), .clkout1(hclk)
);

wire overlay;

// Controller input
`ifdef CONTROLLER_SNES
controller_snes #(.FREQ(50000000)) joy1_snes (
    .clk(mclk), .resetn(resetn), .buttons(joy1_btns),
    .joy_strb(joy1_strb), .joy_clk(joy1_clk), .joy_data(joy1_data)
);
controller_snes #(.FREQ(50000000)) joy2_snes (
    .clk(mclk), .resetn(resetn), .buttons(joy2_btns),
    .joy_strb(joy2_strb), .joy_clk(joy2_clk), .joy_data(joy2_data)
);
`endif

`ifdef CONTROLLER_DS2
controller_ds2 #(.FREQ(50000000)) joy1_ds2 (
    .clk(mclk), .snes_buttons(joy1_btns),
    .ds_clk(ds_clk), .ds_miso(ds_miso), .ds_mosi(ds_mosi), .ds_cs(ds_cs) 
);
controller_ds2 #(.FREQ(50000000)) joy2_ds2 (
   .clk(mclk), .snes_buttons(joy2_btns),
   .ds_clk(ds_clk2), .ds_miso(ds_miso2), .ds_mosi(ds_mosi2), .ds_cs(ds_cs2) 
);
`endif

wire [14:0] overlay_color;
wire [7:0] overlay_x;
wire [7:0] overlay_y;

monitor2hdmi s2h(
    .clk(mclk), .resetn(resetn), 
    .overlay(overlay), .overlay_x(overlay_x), .overlay_y(overlay_y),
    .overlay_color(overlay_color), 
    .clk_pixel(hclk),.clk_5x_pixel(hclk5),
    .tmds_clk_n(tmds_clk_n), .tmds_clk_p(tmds_clk_p),
    .tmds_d_n(tmds_d_n), .tmds_d_p(tmds_d_p)
);

// IOSys for menu, rom loading...
sys #(.CORE_ID(0)) sys (        // CORE ID 0: Monitor
    .clk(mclk), .hclk(hclk), .resetn(resetn),

    // overlay generated by textdisp
    .overlay(overlay), .overlay_x(overlay_x), .overlay_y(overlay_y), .overlay_color(overlay_color),

    // joystick buttons to be sent to companion MCU
    .joy1(joy1_btns), .joy2(joy2_btns),

    // slave SPI connection to the companion MCU
    .sspi_clk(sspi_clk), .sspi_cs(sspi_cs), .sspi_mosi(sspi_mosi), .sspi_miso(sspi_miso)
);

endmodule
